/*
 * Copyright (c) 2024 Andrew Dona-Couch
 * SPDX-License-Identifier: Apache-2.0
 */

`default_nettype none

module cpu (
    input  wire       clk,
    input  wire       rst_n,

    output wire       spi_mosi,
    output wire       spi_select,
    output wire       spi_clk,
    input  wire       spi_miso,

    input  wire       step,
    output wire       busy,
    output wire       halt,
    output wire       trap,

    input  wire [7:0] data_in,
    output wire [7:0] data_out
);

  reg [15:0] pc;
  reg [15:0] inst;
  reg [15:0] accum;
  reg [15:0] bside;

  localparam INST_NOP = 0;
  localparam INST_LOAD_IMM = 1;

  wire executing_ram_inst = inst == INST_LOAD_IMM;

  reg [8:0] state;

  localparam ST_INIT = 0;
  localparam ST_HALT = 1;
  localparam ST_TRAP = 2;
  localparam ST_LOAD_INST0 = 3;
  localparam ST_LOAD_INST1 = 4;
  localparam ST_INST_EXEC0 = 5;
  localparam ST_INST_EXEC1 = 6;

  assign busy = state != ST_INIT & state != ST_HALT & state != ST_TRAP;
  assign halt = state == ST_HALT;
  assign trap = state == ST_TRAP;

  assign data_out = data_in;

  wire [15:0] ram_addr = state == ST_LOAD_INST0 ? pc :
    (state == ST_INST_EXEC0 & inst == INST_LOAD_IMM) ? pc + 2
    : 0;
  wire ram_start_read = state == ST_LOAD_INST0
    | (state == ST_INST_EXEC0 & inst == INST_LOAD_IMM);
  reg [15:0] ram_data_in;
  reg ram_start_write;
  wire [15:0] ram_data_out;
  wire ram_busy;

  spi_ram_controller #(
    .DATA_WIDTH_BYTES(2),
    .ADDR_BITS(16)
  ) spi_ram (
    .clk(clk),
    .rstn(rst_n),
    .spi_miso(spi_miso),
    .spi_select(spi_select),
    .spi_clk_out(spi_clk),
    .spi_mosi(spi_mosi),
    .addr_in(ram_addr),
    .data_in(ram_data_in),
    .start_read(ram_start_read),
    .start_write(ram_start_write),
    .data_out(ram_data_out),
    .busy(ram_busy)
  );

  always @(posedge clk) begin
    if (!rst_n) begin
      state <= ST_INIT;
      pc <= 0;
      inst <= 0;
      accum <= 0;
      bside <= 0;
      ram_data_in <= 0;
      ram_start_write <= 0;
    end else if (~halt & ~trap) begin
      if (state == ST_INIT) begin
        if (step) begin
          state <= ST_LOAD_INST0;
        end
      end else if (state == ST_LOAD_INST0) begin
        state <= ST_LOAD_INST1;
      end else if (state == ST_LOAD_INST1) begin
        if (!ram_busy) begin
          inst <= ram_data_out;
          state <= ST_INST_EXEC0;
        end
      end else if (state == ST_INST_EXEC0) begin
        case (inst)
          INST_NOP: state <= ST_INIT;
          INST_LOAD_IMM: state <= ST_INST_EXEC1;
          default: state <= ST_TRAP;
        endcase
      end else if (state == ST_INST_EXEC1) begin
        if (executing_ram_inst & !ram_busy) begin
          if (inst == INST_LOAD_IMM) begin
            accum <= ram_data_out;
            pc <= pc + 4;
            state <= ST_INIT;
          end
        end
      end
    end
  end

endmodule
